// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
g3SekokMivW2HDRnIkLWxWwv4VHDRrKMTq7I+wSTh0k/67jjnGZhqby/WO23WL/hWD/hZEuJWmcr
D0wUbfiFY+KhmTDez8acXPhzdM7X8ocSmAdQNcdmeVa+SOWu5o4UHAcvYY5+4c40Al5pdrcNyWy0
pz2hnidchXlpPeURzJ2oAisWKZIDhVG5o28oI8SeBljLlghCa+bjouHO78PRWHi5RXO4N3tOXQgX
fM8Fbci/RAmjxjfVLiC2ZyDVeihDSKd4b7+zNkjHmAmLwV/CRilAxKxasRtHtIljMOib+XeJzcUK
KUYvmwvygUa9mmeVYUi2lGgVgMSb3BtbPlYE8A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
bWqzILCi1RtazA9z6vXH3zTjMG88S0OPtX4whhX4bV/0ag8PXVs/UmresjS/8E9UAqIbz6XIDboO
VV+R83PenTH6bN4aMZPHTYojvx6Og6LZCslGBW/HXt9fuS5pd/dMzfLNtyJsDBQuEwZXqmj61+u/
+DRcqzmT7Z1o+Gi1sTkWONRP0M2ggabiUQaczy5SvHzk0XhcXkq9TCbmMy4Zot5uw0xbFws/Jhtw
zO8uEAkYjVsbA/APaarkBRrYwSx3uBk7FhqBwwR6BkKz+JukCb8cPsAAKfAo/r11YYlDYrrU204D
IY1DFvr0s3CJhuIigPRcwPVo8KCDI3M7SV6pKMF+T7PSF/CRk8x5FA9ucQGMT3rnA3UNcFrmFSrl
YlcVKWyWxN0KacJIvK4Y+aiH4OPhU59VsKsYrjpTMqzp4zK7d0AnB5Xzls+PPrpyduVpZjG3HYEj
Eadi20HwDUPy956O5nvnIKbgYrya2T8dp6ktXDleSiHE/sKOt06t1S/RlGYZl4f7/yfMtCMpHnpJ
3ZwDPVw4MHEy0d0Z8XFndW0D8FaaQjOGK3tJzdLibzjbo/6gSxUnnyRXGdaLVWsJfRIR3b7pNwGH
wAzTjsz9Fy81i7ryeGijUAGcy/EUUR3hDkQNPg1OZe8yTEXSRuWhIof/EQvBPBrC6O8tC3ZhUBLM
DHApkpp5nm21Pt83tBF8Kk3ExhVsTIJqXq1yN5mdaHZELBTIlvEDtTGTPqPyqPaJqD22NEqTEu1P
YhJdirv9rhP4cx/G0xwvUkp9IF8yYN+23PedxUhdKr2MWLuJopOohf0dDD7q5WPuwlffAn6laiBC
DQ6VwxIfPN1o2ZaADbFneBNvbQD1kJgiXs1LC4OIIndHC+PPjDpSfYEiRDwq0H/C4tua40GGrmTg
B14hM6CKojtR/FBHMKKXdLuwjfW8JSpu2ycE1ff/wgXw5P/1Fsk7NtYqi6+LvzB209St5p3g1huz
XW3aLDnmM84XHSVa8H/aKhWlhZkn7qwLzCKh3c3tx8OflvBFbrXyTL+4vgaTtY269Sn7rC1c9rcF
rOwwea7nSEG4GDij4q1FOfovigK/a3aQ3h8sd/kohc8obYrCDNaWSBQaZRcD3gfK+HHGvZ+ndTE0
HDS+Z6QKpwOXN96Nxl+hcej0+zoUNv1SWUJ/Nl6JhBGePd9OrVkP9xdKueMRwc/iiGjHiLATr57F
ZU2vmd/JtSnVb/mIVQwiK+f70dKYbf64dvg/pT09Aaj8dYFl1lM8gTjXAQXhCF48Y48Xb79tFhlJ
9MZ4hzmZloCM2xZGHYdqB/1kr63Ml1+jH7IYco88kO+JA8xaguDRk2rQx3n97uP8CVjvvVYyT011
AC2/Sm0x3/ke5vf7rHdqqpLmHyK/sAMNIPjSbBsCoXC3vEplIP5MRoZEYXPCL5QmYWsBHYwhD2fR
qD7ocIKCJZXEMi8beq94S02qqc10R+HzxLKpJtK4+Tx8H/9ogHaARou4PNzjzwXYb2UXuBWfdFjU
CyxXRXb7ekMqqH/Arjmnl2oTbtNkUoxD+0RZeOX8Fo3Broi4kMx6mt0ZJVJLHyhx/BE6qFtH8e02
/PXa8LkhWQnGRLY+2tAB0HXASoEKrUa7jzroknBcZjwZfcJljM8K4TnUANMLTMlx42NuV54fQL7x
fjuVxgEVDBeGRk+fWUUorJTBCDm7hrHfIMYjols/pTs/p31SxkOsUqV/RoujN2oqeJUgaBbpqwJe
iHN99xYIwTEaq1e0JzWGGpzs+/EXLoH3ZMFJL0Hws5YAMmNQW0qouqoQOPI1ZXBnVNLm4I0v6Tor
7GwkDjlSfHH4uCIPsoSOvvf6QZS/Ymlyv/YKShcjckeqXb2rWdTlNw3NDBiOrucjZTM6MULiVlAG
U1bI48ZiAQTCdW/QBrX5RQNzHm/vRoPPekwLlNZ+rD90Q8Wh7W7TLcSa3k81TiN/CutCYlFfcgaL
USnImqB5p+RuGkdXWv0ShCQEvtB5JNyt6DjMVQ+bNIHZMiUzOrupGag//5oSdq54AYxienhBGguU
Q6Y1LLW+YSlicYzCKw5mE2ijSHGvYU5SS6e7rO7LGWoVJ7PsRQe399pZwsvLfCZQs+pUGBdqtvsv
V2fCHF9JzJCIn6rBqm1P8WtJaDAitN2x3xYSCyDVJ3mTx2X8NlIaa8XiehcTtLUIjbS0vi8f22g7
xV8zYpcpoGDiAx34wU+dxTK72T6mg7sN5ucIvAormUUH9+9fVEGmN7lVKhWi4a+xuZLzsdAtmwG3
SqJn9/wKWaorbE3zlilAVoop7rBj31llgGXYOjIXDEVBbpHbNeh8e8c1IAobLrW1Gngek1pD2+Ah
K0Jis1P8NmaH4uaH0fERYP3f7RI87TNozNe1UuIku4KkGQQek8Toutk/TS01iQjFKlHtb09bOqs4
tMbE8E6mnGFzh9uJaGP7yQb4LK3CB10CFm1L6KUFn609l+2nfPM4Pdk1Xe+DpY6UZ0QCsGtllnXk
ouorY7kR3zgBENMxPx6CcwNeQL5maXw8udeQij6FKxAxcMzCYX14svAvoDrstoQ7yi5rKgBtPLGP
EuLgX7yOvkZhzB8nO2Z4iEDHQypQn9XADY9VtkdvMJmTUVH+SF0Ya27GTI3cyErSBvCqUVMrOAyU
AfZdH+S7AIpOB58bYTrLxf4s7OohyhpqPjRQWSy4ta98eChCYoDF2T6kDmc1fibkaV92mYr6jf04
+qmw/BWvx2Xf0X2na5GkfTS1skgJJX37hMHGYYCXscpVTSjy8+qgmOJC6/ICaEzCU6g7ohwomdMr
w+fQkeA/8GTi9jkBsz+nimumrd0yuhnp6tqmJUgUrWdLbwWC9/z7F5Folgo+NVPI+S7xoz/fHqy0
mxaXj+T8Y++qOiasWEhDU1oPJBgXZMgfa2lIzbhxiv8NHjjoKEodQfHPRKzGvTufrVonhDZ6kzPb
YWbmOO0sIvLE2DPMwDWlFDpC7hikULFxRml3B3QhLmpXb2fBkp2NP7ZbLfDa2AT3hMKQvvHZepHb
YMIHYabDaGh4ScS1SPkpwiSX4M4ujFqRtQvjF1N5t06CEb6pSjn7AqK9D6M88eVUR+EaBxJfLxY6
4TusNCn3biQ3LlkJ9MnXtwhG1L8Cf/MEk6Spq8+zmIoikqRIgmrbaWS5atTjpnGAq7DkPY2KrPw+
13T7/XfOim7Z0uxFuL8lXs+mnRXBQuJW5U7s7cecumOY4aZEevTDqFk6UHbqItXK0qzCY84X7mhA
3G14aUCol3DgdUppkEn5kW7Ruw5VR5f+g+kgNRtgfu8OTHShGeMB1dWkEGI20/2WP6HOqtsgLmtm
f9ov6UidmeTkykj/9x56VnIy8OP6pKF3rozi4uP5cta/0jhqRYHhy+KTM7fTad/lp4OLgRV9FJ0b
KzMyT7bw/F7sA1FGxp1D9n4F1v8M2LXpDPftopfkXOxgU9h38NNeSpcwV9+igiiz2s+QRMQTU8eR
A3yGD3c9O77VBM9UhXlopps+Leviy9y5S36ztKNwtIB+4ia/oHSKqzZ2T9A+NYJsFiWK7ywzL6sA
fbXlK4InUSAJkl2+MWJqwZrnJrvehnkLEb9tkuCRYd3BeuKMJwQ36iECGje6Y8k/SQQtNfqqyZvo
4OSjv2w1/lyE3l8bw85c8mXXLGRbthAVeTdMTa/mJQ58OVR2NjZqUdXuYZnmRR/LyR7oSU/L90G7
ZPMq95teFuXpb80iGESYHhc7RyNogSLwJOyXDRyrLtylZA5jvLxlmzLg1V1HqjE0OBbaOrN+JxTD
3gbnkBF8fg+PHrcc4xDTirZ2nKgz/qKbGpNkJ1AzwYWGJG0CofqS1+8J5yFhCWpgLrEKAcpzWCtq
N7vsxOWWUDOE0p1bIH/dpZ5jLWmaRBbNwATx8cPwhKdl6tTOadITSHpFh640WBNqEYDKXcOUWwVj
Jp1qOpnPs8vYhHpPxVU083fHpHPLzvQTjjCiyHXuRKN7Az48B8EhXZu59ViE87utSbMjaIMqaudn
a0+Orpv+BleU6FlRBV5YseUPPj67xuteMshp1k+xhE2ScFpoTc4X2AQ3bIvSKS7FX97XObiz7fue
SMC7v6cjUs3FbiEX7c/hIWtVyfO6UORBVIM+9pEfQnxB5X37sD1FB0j1hq3SBKrci0D58BpjWv/H
dkP7iRVrG1l093Y9XlIASmNAwYcdUr3vqQDS6ebMuQaf/Brqx89y4gYLEdqAu87CkLAI+Raof0g0
1L7JpoTF2hZKgvQLpdrwOjxeYrhrpENdEtrX0CEPohsFwJac+N6paDCft7S3FLlrXWZDieKcFRWX
C9Hl9r5l3jdDGYYm+4q7KPvMy5OFp2GOTY9ovVMLEp+M6WfDrxdtiHDqH2DT6Zs1MHP4IW3Z7A0r
G4lEZHn74emaEaE6l5xkntF1slzAaMwIBYnFGP8WQKUQqZ8RIThQN9AJt8AINnbjDc+vuQ+FR/lE
nkef/4yBXuREoECanGvcqS3FEL/yMiwKbRKQswg+DZOx9OsO0LY2G53jHNFC7Neqk7ljvZ2Jmv3k
+AMSCdlUGYzdIK1gDGioNwYk3bevXoMhUXfS58J+kdCUlajP5ne//s9d/JZvMNzwi3BaG/2gyywh
ULZrd40U/ffBCNkGf1O95Rnf/W8spKaDBXQyK2L863dO7v2+3ET+DoHENBWhOgUedbKpBjjVVuYx
CqTF0BOmecATGSDlcR8R14xBne+paFUZKvm7uLll7utkC2zui8finiaBJZB2c2IstTO1hVsu511M
ts6YzxCn/Hv3ACUheMg67y67K1/FaGbrDBUB1OEshWaw3L3g0GZduMra78xUHF1DcXyslFTX4jWk
ZEGDSOO29fIIh6edDz56RhvWzPAqGCI5arnB8JOUxW8bu7VBuhq4oz73Gm7PD6MJbhdOZQoJND4k
3T4xI0P9usiKfOCkxk8qXi5/C9cDfxgL0uw0k+WT9TspWInTbzlhnfJ0TcwXbl4X4w6OqdMxIXC9
l3SODXKSb5ESOcFJRjhBPp7XwREw2Pv1+2ANgCSEsXmxzwjKmr+6zwRQjZA9z3gT0cniYu+d+qaR
ySDU/LAReTpl26VvuEoG9KwziSeKn728Vqtx6tLvv93WDPfIAYdpXjp/kl8s9fDf2mk9D79BEdgu
FWYnfa39C+EpJRsejrodvt+WN/XTLWFxml7PbOrsViiZrjHXcMj7fxC6NBLXNrQ/s2hajv+mRGJB
uaobbstA+HFkFxJlsX+X8idwSMYJXcJ1kmyq6S69iw4Wl2cVZcVLiBUQcah+lugHgJDkEOYXx4co
1E9gbAfDLUbdMy5v1JmxkSuMiDR5izQbNEPLzVr4W9vp+DSxClrXOjukZR2+AJjv38wb37L8s8+u
ODQfV5Ffch1SWRf9xg1aRk8+e7UZYGypztdJXwBxCnaTAfwEhs5UpHRmEH6xtJcRdqI2Q/2JptHK
q2NJhaSfkrUX93g7Un60WvuipVIgkFRHzimXLawdJADaYmIGTHGSbY32p4nOLaEvY34/XC6sF4k4
T7KMAKnIz+iZPjnb/ojeaRK5omZp+PgQGl9vwpKFq5ABpVMEIhTNZU2S6dFA+zeAmi9BQFNwP2Ic
DO2Lv4OxSzGbb6nzZStsAbi0qzq8DyczjliREopANf7h1y7Dw1EOnn+qLeTI1WM7NQoBHkHTeSzH
ItH4g41I+tsbbw7bn5HtGVWApQWmlcHSBp70BbxIZmIdXBbtcy1ogF4q+a+y96Y886sxv7DlEtGX
uiHIptVnY2Ueun1B8ddtmMO5o8e+/OtMS5Jvoz6JpmidaSTrIocYneYZtGZWggo0YNggk1H4eRnE
6opoQeGgRH0yB36UbiwLkcTqBaUUDL4XXKTgscUV0U5KU5zd7wI4obCEo/X8MKuRcoXukosdFv5L
nbMzBYwsNyBC7fOM7MuPgf1jWo2hWy1fxVGq5z5Ps5VV/cCLnmABIyBZHtXJTN2uwyzrWHPkWvxU
UBtiXkh+v8sFx7bTHQEf8Km+OzXdH4/gMsqtxJtkpSXQXXxLdhioJ0NJyuA5mz4ilVqay+D35mzL
2bXu3UA2sq/ESCZUICVxSTI4LnIyhC+yI2lCNl7Xscdt92cwPxRTFgPuGiVKtQypont7Jk8QAYN6
C0b6Ll95+R15qmYmqzPTfBPf1LcNzFV43w2EzSsbMQ8KKtlm97g9tFpYDaWjYtiHloli7n0Llnwy
HBS9/v2MFCaElIkJY7YnxTc+vb5MCp4REjMIk0BOk8KE5pHnvfBc3GpiPwJn/4Gk4JvIFn5Mn5u/
MFnRMPG/JOSG4bDHmPPgD+TKPMQcGn+otcqq9kRk+5UWDTrzvvM7R8SYwapXYxd2DJnAUNZfS7xI
IJMskmi4iR6SS5/UMj6EuEkeFHXy4iKU5mOyskIgmlzV/Z0itkz5H3Y1z9tw3TWPqvpkkFGbsVe4
d1d1pG5/1PPXMQZc6OAwDQ2nA3N2CvOZ1v+0tWvE1xzpofAYxlxG1rSgl80nyFs6my6V7NZ/PDwo
3V2Lv8z1r/AVROnQcoTwNWdQr95nrufkMg6rBB7v8G6p1xnhl5kwZbY1NNtC5RhhmdkYWqeSQSsK
XN3zbgMZhXQIzjiUKPaA9ACRpFOpKy8uTF2vlpMWYFz/klJ8fua8HQXInoLTkvxghkCyRNlZKChl
Bp236oK6iXzzFLHZ7efh7PBhqb77vXTODZwpJX6I/jgmh+cESFrqmvOTXsTllYqIoWhabUTaTUTE
oM5rg9KJfoViXpVLpC080zU7H6s6kK8Mj0LjvAur20b/xfUJXGJSKxLWZMNwKm4MRPoytWdAKdu4
7YNnWkZT51zl81jub47P6JLdHSRG5F7Fro8+PxKt4EJ/7J3vEb7m820U97P3u8Evj3qBGFH7S80q
rT/Hnh5o+lZlmhQQBLe6q8nA8XWDxw8jGs/x2itUMK4CseB2/FWyjuzd9KPOSPsDf9Or8GU1tRMz
TINja5a3bGLAlyFID8UAKEnSob04zQXpd/vuaTInvWdhKrLrEjJkmkQSzllbnhGyZEMmBVv3nNoV
OapkqXSfLYff3zGq4Itbu8pQM9+Z7XBaZcivDilQ30JiExCS/OsCfJxIIwwGxIMjAcd0Y3xHIMLo
8z8oRpL2okreytvFLLtGyHsxX5ZNzFDZGZJkcS1e6PwYkaTmlz9H3WEghMH8uzQFQDfUuee07XnB
ZNsuHzjFK8zDcM72+6AR9xgaTCeT5YRWH6Zq/eHTLFXqBph5cvlIRNpPmYlxGdK2oOKp5JPcyXJY
1y/VKAPs7sNTEir6+L9A7Tq9hsJ/Z3dTKUXMwPZj/j9Ga5LkRNncQO+V7ve6SA5/tbFH49NDkjzI
SabRq3s4MhA0Mrs2q2hKJDpPyfRpFEpvOauaWFgQY9EvuMEuU19TMnHRreeF7y/CSzjkaTLu1GPt
7VENkjrP7zR/WyR+HaOqZM1Kj6mYYqjeDn5SjvdlSCDBXzgtSm0yMHrmaTJhEsjiM8tvHRsesAcj
6BVLnZJB+pwKmA0DtTZSFtHszkb9jVq+aXRglq7GD049fQADgAqu65ssPicLp/aNfX598pl7Luwr
gLb4aTdpaczRPzaUuOdupeCJYSoMnceL7COe4Mxd/Y9mBDZeyWi7wQGEnvAxDCAltXKNRyK69k3r
a36CreCh9zKQKBZpZJXcqWCY0eG3r5sDmTlHXhsf6iNeMW/D1OnYtbis7Kf2uXWILWvod92Q3poB
vnjAiSLbOiuunhV8Y6VdOjR8bYwtzeGyG6stf1MCxIjEpfgCcPUP/fHmTMLFD3MTVzf+l0acqGh/
TX5Ro2p78QhBlH34pDEJJWaZB72EOXDlyqp1JYSZiphVArQqZeZayMPg+1BsjC28w8xcaQvenWSl
EuLK8O505boWPxnG9Ek4GhYov1SdWdx0D+lParLkuYCJmT/Z2mluGrHcRRUDto1LhogRsEC1bLoJ
Q6juq/eRgJRWYyte7KhUOqCWnK1pv/R0I3Ax4GMcjLW9lFtuN+NtsQaGQAcU1mChXoa1yqv0Ovpi
IsMgikqonWIusOg75grMV3WfnrdGuSse4W8xyk+3UV8Jx73NbgKGLbgJSfVFrx6YGFAJY99XSkod
F4cjzl8lM4g5MqYWB/dnkJ7/pZfgs+i0urQSbuELcwfqWfp/iVv0NcJ1WBYg26KS9bsuZSLudCJJ
Neo22IQezFXytADxnrQxDWFaPHl+tnGJinEMiJ1/SafpQQXiR7pSGKn1uhWD8BO8Y1FX/rMufdDT
CUtkb+FCueNJv6pnGssEral+eaqqzL5QFP4vz62FvdS0DAbutyGfRfRW3z04YmYEeYIYr2/aXRIi
hTjouK6zQ8D4FrD753t7vnKu/hkLouf05U9nUhRYbahsWtLaSV7g+75SAWs/31BHLiCjlXMYiU1Q
mwOchve7KMpXqMmCvcXz2C9eT0yfv6ee2+gACjVkXQc6iR0gRgbEPS4Vy1+7ULAKQmZYrEdUqk4R
sUych26Zen47qVlEYxAkw0i/8xxFI77DeTBoG8AAymo5uHEFjw5kFiUsQE5q8OItT7yr2HnfbvVR
VwCPWp1q3dJlw3IuHBI5td4cttoo6a5WqxNTn+rCB9qOvCEMvt1fnGwxvTWA/oUqEAWiQ7Q25mKo
fgSDmjjN/IPpp+YqYgI9KVVxMb3DLivRX1dJQ9GWN/zG6Bn1/cGsaS15ZNfBxRTgsfr9VV6gZ8Pp
61VJrkJk/ttuMGof+hm15IV5IKCWq4X1LL96GQAw+RT4shodVW5GTS3KqjxZ6A5yYK0yqhiRRUX9
J390Gbtm3ZZhHb8GB2oFrSw7qNS+ZtmKS0Aqh6oNVr1Z1uQHfRMc4rSowdji5AFR+JWAk3daaPed
3kM9KyBZxZGACsmWEvBTSlcXy24j4nfq4KPD/bCvK13vPuSJITmUFJ7Blgt7eeK4Ln37IbXmU7xB
ht/jAytSdSQiQ+uf8exBB1Ti10uO8/fPdOn1G6fcH+IOObZG8i8k/MnVyLq06f7kP9wAyyNT1aGW
9X1i3ThqQBdOpG3ZAgIbkBoOx7B5UkDAi2qvqviAQ0wXv745Q7j+hX2xDgZ90sMnnqrS1zyg0NlX
SlQVtetPpf2szJhUBJXnUaAp7DdItr9mzdufYazndh+MQVjlIPLK5SkCPnepQWJDYSPjdAAPGDXD
2890P0kX4Kl1qG8AMqQGn781nFP5jEGh+43XC61BZjaoyHcV3x1Ef44hT75MbgB1biqOxt4+dPQH
8Lc7YUQSu2bFCqTC79d3EJPxMfYHgN9nn/8iIDZbo11vIbd94019kmhtJZmUaDpDnsWFI5/GkIye
9HSsiffUcv1beSkRN5Ve8AzaNhzW7YRzIHJoQTigDaGMh5fseNQb8qGod39xIAWLgwVNi9vabd6T
fBi1fbVAABQMHRLkb6JSqA27rTlz6/l9SavhATNbBGHdi6bQSkjH9O3Ku7eYbKhNXkOeKmCb+Pc3
UKcX/Ttr5NOb/BOvetyobbZQqpez5cx3p9FCRagQJqfw6SH+Z8gn/QhSWT/tAq79VAyCFh3aLzuc
kdEZCHNTYYmyc2VXGLGa9Av+n09PZu3HSTQ+efQipoXUx9DJJzlwNc/vQLRum+ZKxXDgqmKvZqcE
uerJVQjht7s/YEJv2xDrHNPXR9xRhY+KC465V3yqMbwGoE0aroNsZykI0EQF1xzc2vnszozwZRJn
kz3b+H8dAbI/2PvZh4IGWYMOt/RNPisWBCyzGWyY1n+Ny1DpW51Oty0ZFTf2/eB/U8Be0sy7uCSf
KLWVHcPgf35E9uOeCH0hw91yyKHM1OCrpJb9/pCmvrjQcWQcGOqoTYjn8JctfxvGIcnJlmG+eEKZ
8M35jJsAP/rmCnaSX3J2SmqRM2D83FUgsrtchkNmjWsiZ8SnEcyA44PTFdJCqgi8crXWtT5QQeOH
qadYCdQPHxiXsLtslRi0Fh6C8eGUoRZjgtSPz20tVWtyWIPiCqLgLp5aQrshTdUrnHv3fHmNqBtf
6FUBuTyQ4X4GNrqOkHyvWLn3JyZTrOs/OZagO3PmGTBdtTPMW+lL4TZG8K9P+FSdacFgJ0hv1VDF
AvUZzL+gjmswGz1gfidIxQEz/eKH0oDKFzNcSJor3VAcWH3ANu2hdRvWEaUHFpWE2t2uOiSSeutX
xb337F2uYVMbcaqewSTnR9Zalnl2j5nh3KdJyRVyAWM9G8Zm8UJoAG16O+59Gig6RrBumu1ZsBHE
hLerHT+4T2Sz5JeWbCxINu38gTEqunKduD7hG4Mf3i98y42zSgY4SbBF+OiAn0YndlsO4EjaEyi/
AfvTHupfdwFhn4cerinI6FrjRElS6pSX4d4Gf93zCZCHlMYY0tBk9DVNjM6xqwkFrn+e+62kgXe3
poQKZI2jL+SfG6+U2SCuSgiEATRsvnjTMT3r2eK7vdGsaWJg6Lf03tSSaDwMEr2C2d528uU7XH5v
fP/bLa6bzvA4dOS8NG5P2jdo7rglVppcc8RFxkzmYTW1/fAuuniWh0iQeo0EOO3K1LWpWwi866+5
miYUsQPtjW+nFKEeF8przBdqinYoCFzJVN3zujFD5fRbKtpF47VQCpSWcHPMZ/0pWgz7AVWcyMNl
OigzDUKC3ldzIhs0x1Me0J5OwJXKv0TB+658PbIsjdL8kYe7WIRW158Whu9pwzwycEjzVag317lN
N3oBNqel1VAF2W6M373c7Sg8j2uVpSugCSkj61fgDBS3UbFt72+zRDBki9szpaJLYrurhICu4Hbb
bHBU8ECXrUaz2Ckev9vSTcAf+TdYQui7AjDCYZ2WRQ/xhmZiy2Vz+GGsTLmI+WWTA8+QIyjpo4b9
ewVJ24BU14UY1deJtGK9whTzU8VRpMpUeT/JZ1YKl+71DADkrGvvfh9UXO4QXKGltlRbgp26GGf8
+ae7LWaRRgCl+MZI91GZdYYhbknBBmgdWBCz+Ce07R2K1ymx8wAuh3lILtwXuvJ8zZIh8UolM7s5
Jk05Y0+aVq1uDTWwv3bMlKz+jkO8/yIjf4FQSqTHkKfnIkGOyBqtrRQr+jQv8XVQPWoV04ZgFOec
rMRQNDccWOIWzcSqiDARJa2xx9XK+CpIpZzGkrrX0nFiTD1LwgZSOHAO5cVDAVMbMCTE+rsCTmn2
gamIQeMJ3iogSjXFhCLlniEqLdGSuMI0zPHCiXTB4T9cQvZLU8j0N1bvQbdTVVR+PgPeFjEZ9OY8
ZY9JE0SVEJE5VIU1MOWy8tQk2vaDdfDB3FWYvmYOsIzlNRIxKDUcCrI8otbTxSMAcTvyAkoiSF24
59YdxuESNPdCsFgGJARw4j2KG6lPUK4N7wm96h2bdWunETzEqMxwQRxFVtLjgpGi4b+8czeoR/N9
OKNBhexMqQzo8l0SkMwH4SakN1mFRJSxorc+XXFOkaG8WIPJNIwJpcHGbJUS91NCIJPDrlj7haek
JgS5oDyhowDTXy6WHHKxW7Sp3p/fZJZVhHZoxO04PoJ/yqh8nqYsobkDO2uvLGfJOStKNd0uPy3q
ZJKrD28RMzdcJff7i1ABIte/E16U7JPT57ZS2+lznFKS+8YBEbbVjDIwRcnuwqkvqOpGQvQlVjBV
aqDQpsy2WstBfmQMIQGP68PFIf+mxtfvXYns3+qLjXO4vOw8U4rkIkiKK3dJai2g4qJmfjxs3lBC
RSCBDrluOwjEF6OAxx2eToxPl0GYGLp8ir3rESHLVMXAa0mtSF45fXEM7WSncihL18qvgUIc6fFR
+/q7gCCEWtHrRBqx3NH/D8MyjSG0viacH8WHyQuxF0CwztPAbf/3mFv3K0xy8nZZr6R3RHONHB3T
/H5C2hvsAtVhHgp0PLsRbiKCDjS4H+fmcslUTxDHwY7ZTJjT/cwMiO6221/j1yPW3/kBAWTxoAym
m0a5ZefGQdisdeJ/9F2/GvyaREeKGGadsf9gTLFCdgA83/7D7Vsg/NvF6FWIUcNY13VRBxOZ5jEi
Erxli8rnC8OMdJBXXJl34dfXMsT1xTY1YBQvdbgZFtxa0KXF6Um47tMSGecLDlGv8l9kw00MiyIU
NKrHVQQusDBk66gCpSAQELZAAvTi03k4w4U5ukGc4NkmXRQW4X/+rEjQrhx8C3Eaffiqc4s6xGnf
77N8IHqyGwjIcXWcMc5ZFgqXfftaEHvLgdyCyGopwTlXh+udGUT7LrwM22c8s+t0W7zhe5Zy1r8z
6S1Ds7e9mRxRWCIBfzTerNkw5iEzeRqwKpvPX6jceV7NG7qLczB3XUTZ1kwkgql5CXeLIkaY2LAW
otD7NueZyvxwyY1BQRO/zRezEgfgvEwkJgGwF0KnNYkbmrmlQq85elnUooY9K+gPh/BXr5Ujtp3o
A17rdwUi99NdhY6C6q0/anA2RD+PuA/ne6anAN/4Xb7+Aed+Qv1TpWWsV1DhJoV3UdSHUX/x4v+S
vwloHHca66jXYZqHFuP5ElaMTetteI85tueb2h0uv6GQnKdgVIyZah3oDAOV9uG8hctqphE0wApy
PTugOhDiub7m09279bsKnQOFsQRqXL46in1G70CyVso+neM8BRuxb/cD5+ViHNihE4tF9C4cL2ny
omfx4ZVZ7dYnwa47ZEVoc6p8fToAsT4zxKCYnhekNqgwgIeaRAmJIW/rb/LzHodCR3aRiBjlQa+G
a2yFYq4gqvmiLe/8GhnEe9/jPOAJKd05JhpO0sA5Lr19OCOZo3XhVEU04/OUmcsYxiJ6NtM4pEt6
vIBfgEDYjLsc+3kYAxYnA5HIvKkAD11xmMxK+rmZUB04tP9xfsvxJj5fDlkeaZF9VgyGinlX0AVp
hQdVSpPrpsj8pkmgavFrefbF7S45SxCppVGZw0sUFuzrZNy7Lu4bAIKey07icRQAz2RZ5VqxOP+K
9gBlvOIQYXHC6T8+cMpuaX5bnLH2AVFKkdEYuqx8faeR7L/8G9wM1NtTplCZIdObCxmhc03RQ/Pj
IgHSCjCzNdAdsaP46iJLfyaN/53YbcqT7WcDubY0aF/0T6Y7eg5dbpBSXwIeMdqYi0hSTy+oiEdQ
FPbatZIk83zF3LJfULd68Ep3C0ktxj6UPMd2/HDi4OPATUJ1cieTD86s71iQgCxV6M47ZOi0Lxdr
fa22wDrIZMVJb9MAHb1TjtWasTPUEDzfXLvwBpEkhPIgVUMXcyDISAtByNLI6xxjdCcncxcK3oJW
kGZEDeDwm6j5AdG/CYzYcpuynY1DMPSsD1p0DhrZyp5vGr59Fu0FzzmeAKgyBgvxsbuYiM9ho+Qi
xbLUl39LhXGh6oUUbf5QeFM4cUW5y8psS6hwrjfOCfUh2lGT/nlGTFJ3HpWPCunW9dKnCFiq6xcf
gD98HsY9VzKGA58bxC6B+gmhC0M8nzt1SrWOBR414wTkDBA6hI4a5dbq8Ajk4yRN9axJXac0K3wu
uuYnqbMi3ofCvsjv03xHIJHbwBYObPkOR0dgL28b4gQ6iKF+2DB9MZHKpBldk55tjPDHXFA1KzNR
+5VX2o6z6ugYkehXNqqCNStvOr0sWutXjgnxKYoA+8pip2xQBrewdBXyU+DMB3bZfw1kCwtLFBRc
P9UwdxpeJ1pJhUqVLuruqcFA+mcwJXIRZ4HAzNoO4iIC0vLjHw+GsU4sXXG3NYfx7jF6EcL26MPx
uRzpbgzAyzjbDMPTg69m3KGjW9F4w2LypJhhgrSjV2Qz8RuERw5d9QSgSmyrPEd/UQYwuz+heoAy
WXb3T41rVxgAL0rDz0xLLWM6RN4RgNRacVyhZCIA2gIQgQkGKiTsikmPTbcStpK9/TR9N1lOkpy+
Mk0HKNUC7KKqrZith3AOYwzZ06f8XZha/onwvemuQjHeSmYaQN8c/d1FH6LUH22e2HMoBthgNmC/
9neDYHSy09RY2gCcX17Hlcpd/6z814+e2CB/jz9DPa4CxXBtkP5obT2P9EMOYGqm/oRXQRM+jTg4
DbJFGhAVhM9lehroAjEFLkbqHKIl9n479kOe9PeXJdRBxgWbbpBI1xgLcUvTla6CubV6fNJKQddK
qQMh58zgvW+Fmescwns0JMOYD3oOUlAWkJdHuY9p5gRltUtEPAOl+8WjlrWsxofIA1TjYa5y6D+X
vIvXrdIkVUo44mdCg19LUvFwywRHOJxgts1l39/d83rIsn4D8cBdGQiThPnVku6fxDCroyy+71V+
ycdUMbkzt5ckQlBGs+I4B/cjKBVNLgwWSRZz/e5LctxY4uM4O06mboT0dpirWTSksNqh/FgEhlqs
fK1hO/V+x8JluPExgeEBAtqVjICZ5fKBJdIPjMvodDy6JA3E0PdLH4dxUiOg9ZT938zB/L38162O
Z62Gzsw2hFZzQvAMyBODWPZSUo+dzxqmg57ciiAEa8V7TtUl6IsMr6AuoFwpKrtizWF4ytK4j7IA
ZnMbCTe3Hf9QdRjB532lThSnskU3NRkff5pmcItC8Hrl7edRbtnNEoGAYtrVyghDwnqmNgLgKHio
ki112qDAwgmbcFbjd9F7HZQ5pVuh7tj+oMrgfTOZK8pdI/KP8watkrTDjnhWesCPnT64Dd7Ii6Ny
+j/rIR2mIN3ncJIUuv4y9bNwLp4i9nPMgqoj8c19DRbRZhZK295A2u5gjV0Vb6/JxWKx0/A+KEGg
gq3UpSvwdHz0Ew/cpmWIG11i3LunvOVLvb8ldujWs7cNRpTjBHupFa14WiPT5OQjU8xRcD3+bDZQ
kL5kbpJ5HeY0B35tirSJnj7HELYnPLOg2gXFfCAQh0VFDXY5KdZW1MXUoWAFURBc9sen5blxiDpH
SGJn/n2yxy+YtVM5RapKh3f8kdNKKEkabLB8O7eWTG3N9xgf6xDcjIRSN1CLX+OujM1usqgoAz+o
YZJv/2kA6yS1kvZIixbherwYhctX3wQnp797Ne6krMMQBLC1f2njnYtpvwJnegRc4YiNhgMB10sW
Qs37h7mTh4DaVTsrZNBijmnh7suN6dYDaGhO5TEn3Y3i4DkptDKL+01b1OaSK+MWj2aZajzpxKRg
yO42YYrIgQ2npxulI+mQlsWVDd4rLGr6hZ0w6lVIq7A7dRNCL0wsKnWmNI2oEKvUlTsEUNBLw7uZ
QuXpHAt818dJpJLBfICYUx7zo3rVX3Y9b2b8A3aggFQGPD/kAGqNIcaE3KCi9uWZshrTeYwb5sos
Q8nly/N0MGB7mh9fYDYc2s9v5/HMH7pYCKHhWRRwdoJwKBcuPVzGmJdZ2/3GAtqUtJDvRt0rPU7v
Phl3JWugHYX5zCWzO69xy4UOIazsVM1asHQo1govZTd/bdMQRVKZkFhw5vDuv3HvbTvvEpd8A0AL
wT3jNM6XFc+9XTQSLtLFrO7ZtkN9TVuzVmDbgQ9ASQtZbD3PEMQxyb59M2DaYka80Elt0LcbvGks
xjlvjNwYejMOK7Ny+aGP1ewO/+qkic+p5Nsi421Zb5fcFh6XvKBA+KySoTCJ0UFWyAeuLmUB8pLK
zTjjg9UdADRO7y95yxaQYn8lIlInK6sNY7j8Q48r5p6AeWe9cBLcFoVehS7ZcS95bjDHXoMK+vbm
xJD/yHTjaJTYA7cwqEQDU7ns39cLTSjuLml7uos0eocHFYTPaUPOuThJUMd7mIxLOvGlBv7q0azi
S1fs+dgSDNTcOETaWAygUxmSzeuIJ0xowyZoRWwUrlI8/icPysT/SGSSj4dwOw61a3jdRrH5eB8G
H3rVkDTm+tguSxa2I0DC83jQZ+1DK2hyvYCMqde8yCzT+xvAzy3tNyl9hMBCYoZvctgSFn1iOaiU
wJqxBnnHaoQMyIX7pRdCanMY9WPptKbty/JA6FRZayMSrfojltfDYkYnwy5M5LHpNBSlem9LNMda
e3hqaV4Uf61/SoFsEehCN3in6zTUODYBbcmVFYUDAI0Y71Gu80hdNB+djiJFAWMVMNPkQTCz3cgR
yoqD9rYlaW9zTt9U8O9QRXUHRLWIp4D+hw+6S0L24CZ+ULIDFbXk7f4bp3dcrTw8roE8JWa4aocX
/0avhgHXDPpJzbPWYeU2Qvx0fkzEkCiu009WMD1Gko6VzNBV/ozYApUVkxJNNvZJHmIGNthOBH0K
rlJrOOVf9PyiJy86yH/ceHJlaoDew3d47AnMjLEzW/6IdaVNPh5ZZKaDOmgbGvrwCrfMLtyxujh1
P1LkyIiJm8H/QGo9vPzI/LHaYbQGnUUbAjtYKSUNgX7OGUWxumxVYpmoytsSp5Yy6hYxXFsVqxPV
fjZ0olblUcFZ4R1NpLeI2kKURevQB1J5W4Aet1w9J8KyYNbb5w7lUXszT/Afcl9YuZyIbAs1SkWG
wWdvlz+zrRn5jzm6eAjCvB6RsovA8ngP6ezq963PZrkBIYqLkv71yY+EaWtzyO6vQHk27Vbt7WTp
+mouJwzdWpy6juhj++5Clg5z8WT2OSoIJzdO95oRGJdwC5Sippq8KzeL0G5RaBkEW3sz0c5C7u6L
7sPv5ZhruKzwgav8X5EPsQ31hbWII52qhRk95c2E9C3MAPZyodoi4Hxp4PTEgVkxy0HGh94HVSj8
DrrJ3412bxzBs4RvuEJZiLArQQ2GIEQYcPnZuRU2IfUOssBKk+i2WKJZ7b/Pn7UkjhS10a5jYX2V
DSwjt8uO3iKqiH6ZorjjS5ubYy9SZrVa14ystzQkS89jxLR2fqduPR6szfvJnrUOLsEt0Iz6OrKC
J8/8Q++4KiQdyliWrmWZI3gBi4fXicZ3vVhXi07Y+zkNmoC5IIT7LdyzDp0NPVeT1kxir7uiMFOJ
N3zZZAdIucp5khfhZrJ6Hy3tcDNN4PPE2G1nn9A4PWAJKPtn6uyFXr08UkD0ojKtWWsXkCYepIKL
cQt9zrRwDWRLxJbglcbGD2DBCyFKS6KiNV0aMe10kUGy/sNrjXyiAPehJuwBA/doD7mjYym47Q5m
GmWhII65gCnL7ncEfoe6duhPm9kP1perwSz7u+JHcjOXTv4b7lRz3lFOLo1SCojC6Ys8Ex5nmWBs
98Hu64LZA4/43eWhWxBaC0e+iUjHfkd3q3TrTJ997+7yhREdclwvX9L6FOLFG4YfBP2ggn0fFzrt
gpcTU6yNdu1gMxm3SS9bWf6gnty7SJSfBOKjmq+eY65sRYAdL5PVgPwfFjQN4xqy0qjZXajoHnDL
jI/wGy5dpFOkBXHYkhOkYameOSH/u84P2qa9W82LGE4FZjCARNzWW+Be6V+k2Pli1JyJY+INWOGJ
oVM+NF2sLiZsh8/GZacdqRHT2g+IbTu/A8cHxKENZzA47yVjfm9LO+pehVmoZrkyiV2x9evlCjOE
DuvwUISKyvallBT5POQSUpvTBWeB81PqcjTfBd16Unw5GJIYGXh77THw3Jp8Rb1hWRgB5GcmQaeA
F/U1tcUeTbJHj5XWCq/q659FUMeqB/613uWpm0k0q48Yw0DDDVup4YFAN/gcE5jkopqynHgH0hX4
gKstNwI94PDs2K3rFJtWsgNpjh3x5+EqwvFnpAYM1UdZVBkP5qZFpcPhZkmG7GV9rTmWkkNvmGtp
E+CLzPw/8bkxBFNahNZ3cJb5lcPlaHOBxENMCYt44zAVGqDBxAqGuNmOPrPrlLEtZm6oiSLekTmA
saQvqZlYtY9mgAKubKSEm418j9dBS37PcL9cfc7QhKhONOPXQ0yMggm3+YAmMzbjwxeVIlvMIziv
W8rJe4KhMVTujr4dcZjGAYwBnYYybY+lc81M5RjSxAV5gWJNQAv8fWPxGkEBZuAx1eSNztPqTTvU
FJEqVfjT3V8Cp3qP2UVIotc1+p3xxbsCi9pDwfdT+5sGR4H9gUke4tkvGAgHwkYACr3sx2ketFSV
eioeUJbGk7xfq2pM8llRBnd8b6LXJsorp0/oQsvZbbVZE5Ia2iXRHqKD/XX7WAgQxVzquvdNGcKh
ZR3coFnxbSUK5S3PCKpNUyWodOcYBzddeXhuauGTGKr61yl3ob2HustYjXiYwyjycJxN2oZi7mN2
s7p7hG4IDLwqLzuOpBj52hSapzrnWNLiwzTVqMtHQReuae2rzr37y8SbCS9pF8mNvVwCCJZU8mQY
R5qR/CrN4zxE02sbFNUf57aVgenEQfEp0hQnXnZBRJE86PmsYaAw1K+UNw2CQV3XK+WurPWwdqrN
uRWVgAfk/kiccgBrGfeAs33KESCXmoVJtXHGGZSvaVPOnrfGP3kHFSPddA7C1Sx0Mj4Q1KnetqO1
pi/Ly2bAgy7fuDHP6vrjk3d5mrQueFks+p7TC2d+lzbFhi6vIFWfIiYvpx2feZ8iXy6MILhUXsNC
y5UDA5HKhW6xFkOwxGiN2VQwDis4M12Fe6zkxgy7cu/DB9imSZryowpACiLbWfqalzRuSbAr6/gR
uvnXIvwN93YAZHXL789zsLuT48kuwzhGuyUa1Xlw6bwUkJLJZFe91UeSExS8objWFUdh1g8ZIEQS
yA9NxtdKzosgVlIC1aslcKpGjjcDM1LA6f6qA0PoHsRukkz/9Uhz/mDyTFsB6JZoDqjNE74saGB7
jniUxHlPasXm2nESyzpfuxfUEBz9rYaC3IGciAbhvy/+o2Umy3UMDLx//Kg1B9gvguNUgteyCWyb
SJmCSSg9YtEOLHAdTJgm/EkyYjTizU1NH4mIXEP4eKe0D0jV5qkK/mkPO6Kwgay49r3rGzjmGddl
e7OvqKIP9yCrdE9kXO7ejFYZJhHi0vOV30Ogz8+3Zm3BVUseXwJmZPkgbJJFqZjV8widb0pcszLG
0xGrB8IMs4tlVtk7HrsNZ+h52KRHWWSMTE09QVG88ZpVd0Emv4WIMkXcoaqZmEoQ1ThjFprzJemP
Ar4zUOCRVo49VKlqi9H02CWU3Z4Fyu6lyOrru/AqmkmOHusNJ3FPhh0MAnRDsQPgWt/Nmg++ZXd0
0ZeOVz5D0tQx3ycGbvAwS0cNHIUQkJlHCVZtRhPd9Ke6rzc+neteTPdeZ8KMWcNlEkX7tdBqUqaf
a9+7aIIiIDdRcPK9+7+LsXIFw0l0uPI79mazfpDUUJVAut5aFRkH+0IfJJuoDlV0r/igZ2oTH1Ei
JqwcStNHh6xYxh3RbtrcIte9A8KIMZ5xWE9sUjOjV721H+tq/zFdVJll0w9NdY76pZOlwroGuSDT
oeci7wTjRiio9swtZOGJsfHVCaTefqW7EGXRmHtzv5Ip/QhJhEouwqSzbzgf2NXs2Biy78E6Pc3n
nseYn0JlET9dxtU29LGdYpBXleKUY2cGXdKGCgmnGrYY9rYlb70/5XipyN8lBYnq8ac1UX9r7lvw
Si0mTLAPCIATH8h9pR60WeQ2+kbM1EtmBjDz3ZdnVh6jeexVSOkFYmqfCIIBnfg55d/bKOtCbzL0
9pFyLQTwxaE/tDwjZS8RltgORsgyRfHQjO//B4Y2e5e/qGpraBcgth5DnFF8htCbdx/FurTM5Jvh
3kM180kqy5lOXLwNzA24iVFRy+KZJ+YGaH9SYxBLUc3Xr9j/YaeU2dOtr00X+wq9r1gtshWzQucz
cfrOcSXv0ITugrJ7W+EQEu4GXzCt8bTHhubMKSEJwtdIZ5ltQ7fK1twKXDzaABUsGr6fT+feldko
IUAAzdtra3VWMrF4xfmmcIuWQZaovydw7/LS/dm0xAcH51y+s5XhRUbbDtoJbLODcgYaFh0ocrxE
K5Efxm9+Cv3sABe29j8NJNAlc/oYGydI6jr8BdNYnJwQkYiKdfJH5Dd9mzpPkEJ6EgyX7Lr74cUO
p5/IPSmxUqwb1J61ElMgtmmvH4Mq91Y4MKs+2lxe6pe0YqCGRfOdU6H3gQV9wBagpHUm/80eQCy9
ZT3EScz5LMlEVdmjj28HRrj1jXedFKN9dryaEhSqEqUSFe+OxR1qEqMx7gkdPdLLVMRAd0F5Z/yu
jd8HczjoQ71y8CTwNwfr0vbX7ovKVvkGfFV8Z6rgsHvZtGH/WlzOKykaOrl/qmzZRKjaWfVAzCRi
Ea47qIx41Eue959WtAzLGbl3MpehukxtWw2oGFqyM8VuhMY0ebYZT/+HFXkKlR3XpdonWBPlcC7y
fbffUrsdDQTeD/izAtg3v3oNtsM3qwMbEOyfeB/xzchMj6kCkHxBbsi5F6ycH8h02P/hBCtcEGA6
ARDIKRjOQZ81Wez6HHybQpTQvgDCMjmH6niTY57NSY3GdsNPoA4aGh0/6mkRyLgMCDkzPV246T5J
sYYotjAZsGiFixwcRYhSOToWJcvUHr3uBs9JjMqEdvzaqITX5nYEy1NLqgyqkfHbWadsRdK4fAUB
JB6zWKo1+PhVGdVIhK5SzYdJkDFB2oXUEsW+nRxlbflL2XV2NuPAxkgETGqNk860wWAnLDQE67Mp
s9cKSnGV1CkReS6GgCF570ZEJAZbihnVv2XJuWq9me6z288lh9uuQs7EJZaIHwgvxWGfN25P0SjD
EEI/ic1r95+DMCICBwoSAObLKee18B0Tk1WMsGrfU3XrZlyDtIvz081ZoBY7PUnQRcAkwaRlp/3W
fQKlVyvA/wabzfcjuWC9yllrVvXyMo9r0pmejtvemCd1hroqUSDfcN6KMpXao3pcK8PHtgV58z2w
xZRmWF6iORZaH7HuvYCfgFIdqZyXTsyXD375R0SoWXSRPD5Ud7gI0zfN/+tVoEjO+OL7VzmyzeiM
a0SFf1qVsWb6SOXYNbUaI8wabvnIn5wsAOnPDYrOvk+G8FEfZ2EXa/CJyCs8ElhI6IQdWdqFcCaK
Px/fCDeh6G6YLTGjDkEAFQxeoo0/0lPzJFHsDIZCstjhiVXSCVzSjcWGFFA+x9DPTvz7WZTgEXsF
CKRMJTapDNii7l+Izo1M4VBZF9p+ub8cJUmdbGVtYjoUMhleyZZW/N/SPfvVe13Dt0/O3fvGjgQC
8CB00ud3mhekRy1lv4ACi99kmAAGr3PosRhgAJ0cB1/0knmx3jZYzGpkZeiYjv+0LjrMOAET5skd
FPXqRTwueKDqxPT0oh7msBufl0hXbacknMVbQREsdsc26bpWtI4N2imVxXYY1HgcFLrvGl7o1jOs
PVaBVG72FcYDB++CU7KImz/hsg+HPpptw7XfF5s9xl/CB89SOMciPvA0Imwpfnx3DyxHo8S7iGHl
O8+0Q3rpLOn40WuXqEc9BYSQ0uC3W18t3nOXiiDNQhCHEg0PnT86mmg6ep06I70B0Ems2M2OG8jN
iFd4TWXWPRoWv5hpDwdb93eWfuw3MH4RxaV3pwXiM1pO7ZmxVzCDc1QmERwqMvRpMkpd3h47l5GZ
9k/RJzoyOwoqeiWK/baGqnpfCZNb66KNEyPpxlnXLWTvD0GaYOS2oZpnOwn2BFvBUlOrowea4m/z
HXwhDr8YzsimtJUcqeG8CAkz986a37WxOoISD5ENeP4I36A9D8gGtyvuJHQkIBnIVUdkFGEdPkwm
s5m2Ofb7j1ebH2k7OMjB/Fi6fqNpBoLw1MVtTmZOY6IPdsqQZ1nDdb5J9p0jXVmVwQvdpMq9ywAx
hTuToosdb52ima6S5EdXVi17HCxpgRFlGfq7QgMu6j8+bt4+o45slH6FaKeBEhVAEgoIEBSdvGdS
sl5uEENCWt4D65CgywZqcqLEN7AChN7hlzGeKyasybg+TNAyDZUzJ48ffCjku7LRPlgxPq/WEr5T
qTidKi5/5BqnG7VPNiB96bqGadripZB6RA88tbrUxcsNvWxnIRQi+FdK9b1c9PXSKvN1VwHgQ2T9
L2MTuFi/zBCc3mQyCkMAwRXX/EgPGaG30RciA0zSOuRnSP/x9Q5OnRsoKQlFcixbqwe5kQOwldws
2i/iDBCUVSwXRiEneD+8RG9l0/HL5XH6lKV4ZKKJw0WmpMgrA1a4uZ777LtG1VMxxTL6t/m5XztS
iwgagYN1ZQvTIuFgNQaazJy0GR/ZNI/O+gVYZGqcU7PqfY+RXTWa04oSgjrvvKNbWfXq8aglhJG1
Kw1obOnKvSZ22gi024FW9RS8pq2QYUSGHSWthaediNaPGURTS5XSdxupgABepQPpqf1VIGx1PiGx
RXS1S9CJ6JSUmSqeOiUxFKUMCQWHWJPfNScyv5NoBYC0JejFHCTnqOvRbf3vWpZDIdizF8yzgdc+
SVRqj5WVDG09X/JIwc5WbftVE6fuHsvdYm7UGyn4hJ4l2RHweOdFM3emca1Ih1SvKKD/6GE/eN2p
TrK0dUJVe+RljUMAEQCxzvhzIcf8RUv/V8vPjNvVYBGC2jHomoA8ksRkyglduuWAdciCVFq6vP/5
qTcJMjgyUY2Jly0MjWHC7Cv4oUtiKuX6owJBnm6sWsDfzN5B18JdpGFBB+gTpaucewfZ9sLbx/Kl
siDEccjuXdr9QXBfqyO7brq9cYQNA+X3ctq5RcmGpQe+76ijKBSBdPi+mzDSuln91muiGaGXoTyO
5haw6AkxFwRmzc//bGkXpChZrGaT+B6WogZEpGo/I3S5kcijCeHgbo5sNgKeqhLO++d9KkMXRTDU
J+JcU9oncx0SU6pw48z7Vnus+1/GqUY3DfcegnBZc6Gd5uAFVu/wCvMzyc7JlmshF4t9jxOd1a9w
umw1qmWsXWZ64V82C7Og1bnqJZqZ/iKLJPYkKTYON8/De6C0vZVFq4V7e33oxe72TSbTK7r8J747
O1v9yC5HN/0/lUL2lY0pk8BYS0H5SmAte1adgF8SMPOgyXA3rIOxeipgdb6IyzAMqmScRBhKKxAy
JOPEc7ZoQMuSbo0IzGVdVR94dBfRPdvSvijH+J7Yw/tQLsYo7iuBPQx8HIHT3YRwRo2Fo93HX6HD
7g4jzWz8FWSedZZZLKkVVWxKPYY5vJVvwgadgtTwjIOfG+3wFiljWYAYIPynuJgZes4gLg==
`pragma protect end_protected
