-- lcd.vhd

-- Generated using ACDS version 13.0sp1 232 at 2017.12.31.21:27:04

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity lcd is
	port (
		clk_clk               : in  std_logic                    := '0'; --             clk.clk
		reset_reset_n         : in  std_logic                    := '0'; --           reset.reset_n
		lcd_driver_0_io_io_rs : out std_logic;                           -- lcd_driver_0_io.io_rs
		lcd_driver_0_io_io_rw : out std_logic;                           --                .io_rw
		lcd_driver_0_io_io_en : out std_logic;                           --                .io_en
		lcd_driver_0_io_io_db : out std_logic_vector(7 downto 0)         --                .io_db
	);
end entity lcd;

architecture rtl of lcd is
	component LCD_DRIVER is
		port (
			avmm_address     : in  std_logic_vector(4 downto 0) := (others => 'X'); -- address
			avmm_writedata   : in  std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			avmm_waitrequest : out std_logic;                                       -- waitrequest
			avmm_write       : in  std_logic                    := 'X';             -- write
			rs               : out std_logic;                                       -- io_rs
			rw               : out std_logic;                                       -- io_rw
			en               : out std_logic;                                       -- io_en
			db               : out std_logic_vector(7 downto 0);                    -- io_db
			rstn_sys_clk     : in  std_logic                    := 'X';             -- reset_n
			lcd_clk_250K     : in  std_logic                    := 'X';             -- clk
			sys_clk_50M      : in  std_logic                    := 'X';             -- clk
			rstn_lcd_clk     : in  std_logic                    := 'X'              -- reset_n
		);
	end component LCD_DRIVER;

	component lcd_clk_gen is
		port (
			sys_clk_50M : in  std_logic := 'X'; -- clk
			lcd_clk     : out std_logic;        -- clk
			lcd_rstn    : out std_logic;        -- reset_n
			sys_rstn    : in  std_logic := 'X'  -- reset_n
		);
	end component lcd_clk_gen;

	component lcd_master_0 is
		generic (
			USE_PLI     : integer := 0;
			PLI_PORT    : integer := 50000;
			FIFO_DEPTHS : integer := 2
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			clk_reset_reset      : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			master_read          : out std_logic;                                        -- read
			master_write         : out std_logic;                                        -- write
			master_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			master_reset_reset   : out std_logic                                         -- reset
		);
	end component lcd_master_0;

	component altera_merlin_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(31 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component altera_merlin_master_translator;

	component altera_merlin_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(7 downto 0);                     -- readdata
			uav_writedata            : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(4 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_writedata             : out std_logic_vector(7 downto 0);                     -- writedata
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component altera_merlin_slave_translator;

	component altera_merlin_master_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			av_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			av_write                : in  std_logic                     := 'X';             -- write
			av_read                 : in  std_logic                     := 'X';             -- read
			av_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			av_waitrequest          : out std_logic;                                        -- waitrequest
			av_readdatavalid        : out std_logic;                                        -- readdatavalid
			av_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_lock                 : in  std_logic                     := 'X';             -- lock
			cp_valid                : out std_logic;                                        -- valid
			cp_data                 : out std_logic_vector(98 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_endofpacket          : out std_logic;                                        -- endofpacket
			cp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : in  std_logic                     := 'X';             -- valid
			rp_data                 : in  std_logic_vector(98 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                        -- ready
			av_response             : out std_logic_vector(1 downto 0);                     -- response
			av_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                         -- writeresponsevalid
		);
	end component altera_merlin_master_agent;

	component altera_merlin_slave_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(31 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(0 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(7 downto 0);                     -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(71 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(71 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(72 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(72 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(9 downto 0);                     -- data
			m0_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                        -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component altera_merlin_slave_agent;

	component altera_avalon_sc_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(72 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_data          : out std_logic_vector(72 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component altera_avalon_sc_fifo;

	component lcd_addr_router is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(98 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(98 downto 0);                    -- data
			src_channel        : out std_logic_vector(0 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component lcd_addr_router;

	component lcd_id_router is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(71 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(71 downto 0);                    -- data
			src_channel        : out std_logic_vector(0 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component lcd_id_router;

	component altera_merlin_burst_adapter is
		generic (
			PKT_ADDR_H                : integer := 79;
			PKT_ADDR_L                : integer := 48;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BYTE_CNT_H            : integer := 5;
			PKT_BYTE_CNT_L            : integer := 0;
			PKT_BYTEEN_H              : integer := 83;
			PKT_BYTEEN_L              : integer := 80;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 88;
			PKT_BURST_TYPE_L          : integer := 87;
			PKT_BURSTWRAP_H           : integer := 11;
			PKT_BURSTWRAP_L           : integer := 6;
			PKT_TRANS_COMPRESSED_READ : integer := 14;
			PKT_TRANS_WRITE           : integer := 13;
			PKT_TRANS_READ            : integer := 12;
			OUT_NARROW_SIZE           : integer := 0;
			IN_NARROW_SIZE            : integer := 0;
			OUT_FIXED                 : integer := 0;
			OUT_COMPLETE_WRAP         : integer := 0;
			ST_DATA_W                 : integer := 89;
			ST_CHANNEL_W              : integer := 8;
			OUT_BYTE_CNT_H            : integer := 5;
			OUT_BURSTWRAP_H           : integer := 11;
			COMPRESSED_READ_SUPPORT   : integer := 1;
			BYTEENABLE_SYNTHESIS      : integer := 0;
			PIPE_INPUTS               : integer := 0;
			NO_WRAP_SUPPORT           : integer := 0;
			BURSTWRAP_CONST_MASK      : integer := 0;
			BURSTWRAP_CONST_VALUE     : integer := -1
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			sink0_valid           : in  std_logic                     := 'X';             -- valid
			sink0_data            : in  std_logic_vector(71 downto 0) := (others => 'X'); -- data
			sink0_channel         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- channel
			sink0_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			sink0_ready           : out std_logic;                                        -- ready
			source0_valid         : out std_logic;                                        -- valid
			source0_data          : out std_logic_vector(71 downto 0);                    -- data
			source0_channel       : out std_logic_vector(0 downto 0);                     -- channel
			source0_startofpacket : out std_logic;                                        -- startofpacket
			source0_endofpacket   : out std_logic;                                        -- endofpacket
			source0_ready         : in  std_logic                     := 'X'              -- ready
		);
	end component altera_merlin_burst_adapter;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in1  : in  std_logic := 'X'; -- reset
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component altera_reset_controller;

	component lcd_cmd_xbar_demux is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(98 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(98 downto 0);                    -- data
			src0_channel       : out std_logic_vector(0 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component lcd_cmd_xbar_demux;

	component lcd_width_adapter is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			in_valid             : in  std_logic                     := 'X';             -- valid
			in_channel           : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                     := 'X';             -- endofpacket
			in_ready             : out std_logic;                                        -- ready
			in_data              : in  std_logic_vector(98 downto 0) := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                        -- endofpacket
			out_data             : out std_logic_vector(71 downto 0);                    -- data
			out_channel          : out std_logic_vector(0 downto 0);                     -- channel
			out_valid            : out std_logic;                                        -- valid
			out_ready            : in  std_logic                     := 'X';             -- ready
			out_startofpacket    : out std_logic;                                        -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)  := (others => 'X')  -- data
		);
	end component lcd_width_adapter;

	component lcd_width_adapter_001 is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			in_valid             : in  std_logic                     := 'X';             -- valid
			in_channel           : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                     := 'X';             -- endofpacket
			in_ready             : out std_logic;                                        -- ready
			in_data              : in  std_logic_vector(71 downto 0) := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                        -- endofpacket
			out_data             : out std_logic_vector(98 downto 0);                    -- data
			out_channel          : out std_logic_vector(0 downto 0);                     -- channel
			out_valid            : out std_logic;                                        -- valid
			out_ready            : in  std_logic                     := 'X';             -- ready
			out_startofpacket    : out std_logic;                                        -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)  := (others => 'X')  -- data
		);
	end component lcd_width_adapter_001;

	signal lcd_clk_gen_0_lcd_clk_clk                                                                      : std_logic;                     -- lcd_clk_gen_0:lcd_clk -> LCD_Driver_0:lcd_clk_250K
	signal master_0_master_waitrequest                                                                    : std_logic;                     -- master_0_master_translator:av_waitrequest -> master_0:master_waitrequest
	signal master_0_master_writedata                                                                      : std_logic_vector(31 downto 0); -- master_0:master_writedata -> master_0_master_translator:av_writedata
	signal master_0_master_address                                                                        : std_logic_vector(31 downto 0); -- master_0:master_address -> master_0_master_translator:av_address
	signal master_0_master_write                                                                          : std_logic;                     -- master_0:master_write -> master_0_master_translator:av_write
	signal master_0_master_read                                                                           : std_logic;                     -- master_0:master_read -> master_0_master_translator:av_read
	signal master_0_master_readdata                                                                       : std_logic_vector(31 downto 0); -- master_0_master_translator:av_readdata -> master_0:master_readdata
	signal master_0_master_byteenable                                                                     : std_logic_vector(3 downto 0);  -- master_0:master_byteenable -> master_0_master_translator:av_byteenable
	signal master_0_master_readdatavalid                                                                  : std_logic;                     -- master_0_master_translator:av_readdatavalid -> master_0:master_readdatavalid
	signal lcd_driver_0_avalon_slave_translator_avalon_anti_slave_0_waitrequest                           : std_logic;                     -- LCD_Driver_0:avmm_waitrequest -> LCD_Driver_0_avalon_slave_translator:av_waitrequest
	signal lcd_driver_0_avalon_slave_translator_avalon_anti_slave_0_writedata                             : std_logic_vector(7 downto 0);  -- LCD_Driver_0_avalon_slave_translator:av_writedata -> LCD_Driver_0:avmm_writedata
	signal lcd_driver_0_avalon_slave_translator_avalon_anti_slave_0_address                               : std_logic_vector(4 downto 0);  -- LCD_Driver_0_avalon_slave_translator:av_address -> LCD_Driver_0:avmm_address
	signal lcd_driver_0_avalon_slave_translator_avalon_anti_slave_0_write                                 : std_logic;                     -- LCD_Driver_0_avalon_slave_translator:av_write -> LCD_Driver_0:avmm_write
	signal master_0_master_translator_avalon_universal_master_0_waitrequest                               : std_logic;                     -- master_0_master_translator_avalon_universal_master_0_agent:av_waitrequest -> master_0_master_translator:uav_waitrequest
	signal master_0_master_translator_avalon_universal_master_0_burstcount                                : std_logic_vector(2 downto 0);  -- master_0_master_translator:uav_burstcount -> master_0_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal master_0_master_translator_avalon_universal_master_0_writedata                                 : std_logic_vector(31 downto 0); -- master_0_master_translator:uav_writedata -> master_0_master_translator_avalon_universal_master_0_agent:av_writedata
	signal master_0_master_translator_avalon_universal_master_0_address                                   : std_logic_vector(31 downto 0); -- master_0_master_translator:uav_address -> master_0_master_translator_avalon_universal_master_0_agent:av_address
	signal master_0_master_translator_avalon_universal_master_0_lock                                      : std_logic;                     -- master_0_master_translator:uav_lock -> master_0_master_translator_avalon_universal_master_0_agent:av_lock
	signal master_0_master_translator_avalon_universal_master_0_write                                     : std_logic;                     -- master_0_master_translator:uav_write -> master_0_master_translator_avalon_universal_master_0_agent:av_write
	signal master_0_master_translator_avalon_universal_master_0_read                                      : std_logic;                     -- master_0_master_translator:uav_read -> master_0_master_translator_avalon_universal_master_0_agent:av_read
	signal master_0_master_translator_avalon_universal_master_0_readdata                                  : std_logic_vector(31 downto 0); -- master_0_master_translator_avalon_universal_master_0_agent:av_readdata -> master_0_master_translator:uav_readdata
	signal master_0_master_translator_avalon_universal_master_0_debugaccess                               : std_logic;                     -- master_0_master_translator:uav_debugaccess -> master_0_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal master_0_master_translator_avalon_universal_master_0_byteenable                                : std_logic_vector(3 downto 0);  -- master_0_master_translator:uav_byteenable -> master_0_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal master_0_master_translator_avalon_universal_master_0_readdatavalid                             : std_logic;                     -- master_0_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> master_0_master_translator:uav_readdatavalid
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest             : std_logic;                     -- LCD_Driver_0_avalon_slave_translator:uav_waitrequest -> LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount              : std_logic_vector(0 downto 0);  -- LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> LCD_Driver_0_avalon_slave_translator:uav_burstcount
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata               : std_logic_vector(7 downto 0);  -- LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> LCD_Driver_0_avalon_slave_translator:uav_writedata
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address                 : std_logic_vector(31 downto 0); -- LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_address -> LCD_Driver_0_avalon_slave_translator:uav_address
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write                   : std_logic;                     -- LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_write -> LCD_Driver_0_avalon_slave_translator:uav_write
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock                    : std_logic;                     -- LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_lock -> LCD_Driver_0_avalon_slave_translator:uav_lock
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read                    : std_logic;                     -- LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_read -> LCD_Driver_0_avalon_slave_translator:uav_read
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata                : std_logic_vector(7 downto 0);  -- LCD_Driver_0_avalon_slave_translator:uav_readdata -> LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid           : std_logic;                     -- LCD_Driver_0_avalon_slave_translator:uav_readdatavalid -> LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess             : std_logic;                     -- LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> LCD_Driver_0_avalon_slave_translator:uav_debugaccess
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable              : std_logic_vector(0 downto 0);  -- LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> LCD_Driver_0_avalon_slave_translator:uav_byteenable
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket      : std_logic;                     -- LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid            : std_logic;                     -- LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket    : std_logic;                     -- LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data             : std_logic_vector(72 downto 0); -- LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready            : std_logic;                     -- LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket   : std_logic;                     -- LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid         : std_logic;                     -- LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket : std_logic;                     -- LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data          : std_logic_vector(72 downto 0); -- LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready         : std_logic;                     -- LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid       : std_logic;                     -- LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data        : std_logic_vector(9 downto 0);  -- LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready       : std_logic;                     -- LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal master_0_master_translator_avalon_universal_master_0_agent_cp_endofpacket                      : std_logic;                     -- master_0_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	signal master_0_master_translator_avalon_universal_master_0_agent_cp_valid                            : std_logic;                     -- master_0_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	signal master_0_master_translator_avalon_universal_master_0_agent_cp_startofpacket                    : std_logic;                     -- master_0_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	signal master_0_master_translator_avalon_universal_master_0_agent_cp_data                             : std_logic_vector(98 downto 0); -- master_0_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	signal master_0_master_translator_avalon_universal_master_0_agent_cp_ready                            : std_logic;                     -- addr_router:sink_ready -> master_0_master_translator_avalon_universal_master_0_agent:cp_ready
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket             : std_logic;                     -- LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid                   : std_logic;                     -- LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket           : std_logic;                     -- LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data                    : std_logic_vector(71 downto 0); -- LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	signal lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready                   : std_logic;                     -- id_router:sink_ready -> LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal burst_adapter_source0_endofpacket                                                              : std_logic;                     -- burst_adapter:source0_endofpacket -> LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_source0_valid                                                                    : std_logic;                     -- burst_adapter:source0_valid -> LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_source0_startofpacket                                                            : std_logic;                     -- burst_adapter:source0_startofpacket -> LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_source0_data                                                                     : std_logic_vector(71 downto 0); -- burst_adapter:source0_data -> LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_source0_ready                                                                    : std_logic;                     -- LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	signal burst_adapter_source0_channel                                                                  : std_logic_vector(0 downto 0);  -- burst_adapter:source0_channel -> LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal rst_controller_reset_out_reset                                                                 : std_logic;                     -- rst_controller:reset_out -> [LCD_Driver_0_avalon_slave_translator:reset, LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent:reset, LCD_Driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, burst_adapter:reset, cmd_xbar_demux:reset, id_router:reset, master_0_master_translator:reset, master_0_master_translator_avalon_universal_master_0_agent:reset, rsp_xbar_demux:reset, rst_controller_reset_out_reset:in, width_adapter:reset, width_adapter_001:reset]
	signal rst_controller_001_reset_out_reset                                                             : std_logic;                     -- rst_controller_001:reset_out -> rst_controller_001_reset_out_reset:in
	signal lcd_clk_gen_0_reset_source_reset                                                               : std_logic;                     -- lcd_clk_gen_0:lcd_rstn -> lcd_clk_gen_0_reset_source_reset:in
	signal cmd_xbar_demux_src0_endofpacket                                                                : std_logic;                     -- cmd_xbar_demux:src0_endofpacket -> width_adapter:in_endofpacket
	signal cmd_xbar_demux_src0_valid                                                                      : std_logic;                     -- cmd_xbar_demux:src0_valid -> width_adapter:in_valid
	signal cmd_xbar_demux_src0_startofpacket                                                              : std_logic;                     -- cmd_xbar_demux:src0_startofpacket -> width_adapter:in_startofpacket
	signal cmd_xbar_demux_src0_data                                                                       : std_logic_vector(98 downto 0); -- cmd_xbar_demux:src0_data -> width_adapter:in_data
	signal cmd_xbar_demux_src0_channel                                                                    : std_logic_vector(0 downto 0);  -- cmd_xbar_demux:src0_channel -> width_adapter:in_channel
	signal rsp_xbar_demux_src0_endofpacket                                                                : std_logic;                     -- rsp_xbar_demux:src0_endofpacket -> master_0_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_demux_src0_valid                                                                      : std_logic;                     -- rsp_xbar_demux:src0_valid -> master_0_master_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_demux_src0_startofpacket                                                              : std_logic;                     -- rsp_xbar_demux:src0_startofpacket -> master_0_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_demux_src0_data                                                                       : std_logic_vector(98 downto 0); -- rsp_xbar_demux:src0_data -> master_0_master_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_demux_src0_channel                                                                    : std_logic_vector(0 downto 0);  -- rsp_xbar_demux:src0_channel -> master_0_master_translator_avalon_universal_master_0_agent:rp_channel
	signal addr_router_src_endofpacket                                                                    : std_logic;                     -- addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	signal addr_router_src_valid                                                                          : std_logic;                     -- addr_router:src_valid -> cmd_xbar_demux:sink_valid
	signal addr_router_src_startofpacket                                                                  : std_logic;                     -- addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	signal addr_router_src_data                                                                           : std_logic_vector(98 downto 0); -- addr_router:src_data -> cmd_xbar_demux:sink_data
	signal addr_router_src_channel                                                                        : std_logic_vector(0 downto 0);  -- addr_router:src_channel -> cmd_xbar_demux:sink_channel
	signal addr_router_src_ready                                                                          : std_logic;                     -- cmd_xbar_demux:sink_ready -> addr_router:src_ready
	signal rsp_xbar_demux_src0_ready                                                                      : std_logic;                     -- master_0_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux:src0_ready
	signal cmd_xbar_demux_src0_ready                                                                      : std_logic;                     -- width_adapter:in_ready -> cmd_xbar_demux:src0_ready
	signal width_adapter_src_endofpacket                                                                  : std_logic;                     -- width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	signal width_adapter_src_valid                                                                        : std_logic;                     -- width_adapter:out_valid -> burst_adapter:sink0_valid
	signal width_adapter_src_startofpacket                                                                : std_logic;                     -- width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	signal width_adapter_src_data                                                                         : std_logic_vector(71 downto 0); -- width_adapter:out_data -> burst_adapter:sink0_data
	signal width_adapter_src_ready                                                                        : std_logic;                     -- burst_adapter:sink0_ready -> width_adapter:out_ready
	signal width_adapter_src_channel                                                                      : std_logic_vector(0 downto 0);  -- width_adapter:out_channel -> burst_adapter:sink0_channel
	signal id_router_src_endofpacket                                                                      : std_logic;                     -- id_router:src_endofpacket -> width_adapter_001:in_endofpacket
	signal id_router_src_valid                                                                            : std_logic;                     -- id_router:src_valid -> width_adapter_001:in_valid
	signal id_router_src_startofpacket                                                                    : std_logic;                     -- id_router:src_startofpacket -> width_adapter_001:in_startofpacket
	signal id_router_src_data                                                                             : std_logic_vector(71 downto 0); -- id_router:src_data -> width_adapter_001:in_data
	signal id_router_src_channel                                                                          : std_logic_vector(0 downto 0);  -- id_router:src_channel -> width_adapter_001:in_channel
	signal id_router_src_ready                                                                            : std_logic;                     -- width_adapter_001:in_ready -> id_router:src_ready
	signal width_adapter_001_src_endofpacket                                                              : std_logic;                     -- width_adapter_001:out_endofpacket -> rsp_xbar_demux:sink_endofpacket
	signal width_adapter_001_src_valid                                                                    : std_logic;                     -- width_adapter_001:out_valid -> rsp_xbar_demux:sink_valid
	signal width_adapter_001_src_startofpacket                                                            : std_logic;                     -- width_adapter_001:out_startofpacket -> rsp_xbar_demux:sink_startofpacket
	signal width_adapter_001_src_data                                                                     : std_logic_vector(98 downto 0); -- width_adapter_001:out_data -> rsp_xbar_demux:sink_data
	signal width_adapter_001_src_ready                                                                    : std_logic;                     -- rsp_xbar_demux:sink_ready -> width_adapter_001:out_ready
	signal width_adapter_001_src_channel                                                                  : std_logic_vector(0 downto 0);  -- width_adapter_001:out_channel -> rsp_xbar_demux:sink_channel
	signal reset_reset_n_ports_inv                                                                        : std_logic;                     -- reset_reset_n:inv -> [master_0:clk_reset_reset, rst_controller:reset_in0]
	signal rst_controller_reset_out_reset_ports_inv                                                       : std_logic;                     -- rst_controller_reset_out_reset:inv -> [LCD_Driver_0:rstn_sys_clk, lcd_clk_gen_0:sys_rstn]
	signal rst_controller_001_reset_out_reset_ports_inv                                                   : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> LCD_Driver_0:rstn_lcd_clk
	signal lcd_clk_gen_0_reset_source_reset_ports_inv                                                     : std_logic;                     -- lcd_clk_gen_0_reset_source_reset:inv -> rst_controller_001:reset_in0

begin

	lcd_driver_0 : component LCD_DRIVER
		port map (
			avmm_address     => lcd_driver_0_avalon_slave_translator_avalon_anti_slave_0_address,     -- avalon_slave.address
			avmm_writedata   => lcd_driver_0_avalon_slave_translator_avalon_anti_slave_0_writedata,   --             .writedata
			avmm_waitrequest => lcd_driver_0_avalon_slave_translator_avalon_anti_slave_0_waitrequest, --             .waitrequest
			avmm_write       => lcd_driver_0_avalon_slave_translator_avalon_anti_slave_0_write,       --             .write
			rs               => lcd_driver_0_io_io_rs,                                                --           io.io_rs
			rw               => lcd_driver_0_io_io_rw,                                                --             .io_rw
			en               => lcd_driver_0_io_io_en,                                                --             .io_en
			db               => lcd_driver_0_io_io_db,                                                --             .io_db
			rstn_sys_clk     => rst_controller_reset_out_reset_ports_inv,                             --      reset_n.reset_n
			lcd_clk_250K     => lcd_clk_gen_0_lcd_clk_clk,                                            -- lcd_clk_250k.clk
			sys_clk_50M      => clk_clk,                                                              --  sys_clk_50M.clk
			rstn_lcd_clk     => rst_controller_001_reset_out_reset_ports_inv                          --  reset_n_lcd.reset_n
		);

	lcd_clk_gen_0 : component lcd_clk_gen
		port map (
			sys_clk_50M => clk_clk,                                  --      sys_clk.clk
			lcd_clk     => lcd_clk_gen_0_lcd_clk_clk,                --      lcd_clk.clk
			lcd_rstn    => lcd_clk_gen_0_reset_source_reset,         -- reset_source.reset_n
			sys_rstn    => rst_controller_reset_out_reset_ports_inv  --  reset_n_sys.reset_n
		);

	master_0 : component lcd_master_0
		generic map (
			USE_PLI     => 0,
			PLI_PORT    => 50000,
			FIFO_DEPTHS => 2
		)
		port map (
			clk_clk              => clk_clk,                       --          clk.clk
			clk_reset_reset      => reset_reset_n_ports_inv,       --    clk_reset.reset
			master_address       => master_0_master_address,       --       master.address
			master_readdata      => master_0_master_readdata,      --             .readdata
			master_read          => master_0_master_read,          --             .read
			master_write         => master_0_master_write,         --             .write
			master_writedata     => master_0_master_writedata,     --             .writedata
			master_waitrequest   => master_0_master_waitrequest,   --             .waitrequest
			master_readdatavalid => master_0_master_readdatavalid, --             .readdatavalid
			master_byteenable    => master_0_master_byteenable,    --             .byteenable
			master_reset_reset   => open                           -- master_reset.reset
		);

	master_0_master_translator : component altera_merlin_master_translator
		generic map (
			AV_ADDRESS_W                => 32,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 32,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => clk_clk,                                                            --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                     --                     reset.reset
			uav_address              => master_0_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => master_0_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => master_0_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => master_0_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => master_0_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => master_0_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => master_0_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => master_0_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => master_0_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => master_0_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => master_0_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => master_0_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => master_0_master_waitrequest,                                        --                          .waitrequest
			av_byteenable            => master_0_master_byteenable,                                         --                          .byteenable
			av_read                  => master_0_master_read,                                               --                          .read
			av_readdata              => master_0_master_readdata,                                           --                          .readdata
			av_readdatavalid         => master_0_master_readdatavalid,                                      --                          .readdatavalid
			av_write                 => master_0_master_write,                                              --                          .write
			av_writedata             => master_0_master_writedata,                                          --                          .writedata
			av_burstcount            => "1",                                                                --               (terminated)
			av_beginbursttransfer    => '0',                                                                --               (terminated)
			av_begintransfer         => '0',                                                                --               (terminated)
			av_chipselect            => '0',                                                                --               (terminated)
			av_lock                  => '0',                                                                --               (terminated)
			av_debugaccess           => '0',                                                                --               (terminated)
			uav_clken                => open,                                                               --               (terminated)
			av_clken                 => '1',                                                                --               (terminated)
			uav_response             => "00",                                                               --               (terminated)
			av_response              => open,                                                               --               (terminated)
			uav_writeresponserequest => open,                                                               --               (terminated)
			uav_writeresponsevalid   => '0',                                                                --               (terminated)
			av_writeresponserequest  => '0',                                                                --               (terminated)
			av_writeresponsevalid    => open                                                                --               (terminated)
		);

	lcd_driver_0_avalon_slave_translator : component altera_merlin_slave_translator
		generic map (
			AV_ADDRESS_W                   => 5,
			AV_DATA_W                      => 8,
			UAV_DATA_W                     => 8,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 1,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 1,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 1,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                              --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                       --                    reset.reset
			uav_address              => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => lcd_driver_0_avalon_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => lcd_driver_0_avalon_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_writedata             => lcd_driver_0_avalon_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_waitrequest           => lcd_driver_0_avalon_slave_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_read                  => open,                                                                                 --              (terminated)
			av_readdata              => "10101101",                                                                           --              (terminated)
			av_begintransfer         => open,                                                                                 --              (terminated)
			av_beginbursttransfer    => open,                                                                                 --              (terminated)
			av_burstcount            => open,                                                                                 --              (terminated)
			av_byteenable            => open,                                                                                 --              (terminated)
			av_readdatavalid         => '0',                                                                                  --              (terminated)
			av_writebyteenable       => open,                                                                                 --              (terminated)
			av_lock                  => open,                                                                                 --              (terminated)
			av_chipselect            => open,                                                                                 --              (terminated)
			av_clken                 => open,                                                                                 --              (terminated)
			uav_clken                => '0',                                                                                  --              (terminated)
			av_debugaccess           => open,                                                                                 --              (terminated)
			av_outputenable          => open,                                                                                 --              (terminated)
			uav_response             => open,                                                                                 --              (terminated)
			av_response              => "00",                                                                                 --              (terminated)
			uav_writeresponserequest => '0',                                                                                  --              (terminated)
			uav_writeresponsevalid   => open,                                                                                 --              (terminated)
			av_writeresponserequest  => open,                                                                                 --              (terminated)
			av_writeresponsevalid    => '0'                                                                                   --              (terminated)
		);

	master_0_master_translator_avalon_universal_master_0_agent : component altera_merlin_master_agent
		generic map (
			PKT_PROTECTION_H          => 92,
			PKT_PROTECTION_L          => 90,
			PKT_BEGIN_BURST           => 85,
			PKT_BURSTWRAP_H           => 77,
			PKT_BURSTWRAP_L           => 77,
			PKT_BURST_SIZE_H          => 80,
			PKT_BURST_SIZE_L          => 78,
			PKT_BURST_TYPE_H          => 82,
			PKT_BURST_TYPE_L          => 81,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_TRANS_EXCLUSIVE       => 73,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 87,
			PKT_DEST_ID_H             => 88,
			PKT_DEST_ID_L             => 88,
			PKT_THREAD_ID_H           => 89,
			PKT_THREAD_ID_L           => 89,
			PKT_CACHE_H               => 96,
			PKT_CACHE_L               => 93,
			PKT_DATA_SIDEBAND_H       => 84,
			PKT_DATA_SIDEBAND_L       => 84,
			PKT_QOS_H                 => 86,
			PKT_QOS_L                 => 86,
			PKT_ADDR_SIDEBAND_H       => 83,
			PKT_ADDR_SIDEBAND_L       => 83,
			PKT_RESPONSE_STATUS_H     => 98,
			PKT_RESPONSE_STATUS_L     => 97,
			ST_DATA_W                 => 99,
			ST_CHANNEL_W              => 1,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 0,
			BURSTWRAP_VALUE           => 1,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                     --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			av_address              => master_0_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => master_0_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => master_0_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => master_0_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => master_0_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => master_0_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => master_0_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => master_0_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => master_0_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => master_0_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => master_0_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => master_0_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => master_0_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => master_0_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => master_0_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => master_0_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_demux_src0_valid,                                                   --        rp.valid
			rp_data                 => rsp_xbar_demux_src0_data,                                                    --          .data
			rp_channel              => rsp_xbar_demux_src0_channel,                                                 --          .channel
			rp_startofpacket        => rsp_xbar_demux_src0_startofpacket,                                           --          .startofpacket
			rp_endofpacket          => rsp_xbar_demux_src0_endofpacket,                                             --          .endofpacket
			rp_ready                => rsp_xbar_demux_src0_ready,                                                   --          .ready
			av_response             => open,                                                                        -- (terminated)
			av_writeresponserequest => '0',                                                                         -- (terminated)
			av_writeresponsevalid   => open                                                                         -- (terminated)
		);

	lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 7,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 58,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 8,
			PKT_BYTEEN_L              => 8,
			PKT_ADDR_H                => 40,
			PKT_ADDR_L                => 9,
			PKT_TRANS_COMPRESSED_READ => 41,
			PKT_TRANS_POSTED          => 42,
			PKT_TRANS_WRITE           => 43,
			PKT_TRANS_READ            => 44,
			PKT_TRANS_LOCK            => 45,
			PKT_SRC_ID_H              => 60,
			PKT_SRC_ID_L              => 60,
			PKT_DEST_ID_H             => 61,
			PKT_DEST_ID_L             => 61,
			PKT_BURSTWRAP_H           => 50,
			PKT_BURSTWRAP_L           => 50,
			PKT_BYTE_CNT_H            => 49,
			PKT_BYTE_CNT_L            => 47,
			PKT_PROTECTION_H          => 65,
			PKT_PROTECTION_L          => 63,
			PKT_RESPONSE_STATUS_H     => 71,
			PKT_RESPONSE_STATUS_L     => 70,
			PKT_BURST_SIZE_H          => 53,
			PKT_BURST_SIZE_L          => 51,
			ST_CHANNEL_W              => 1,
			ST_DATA_W                 => 72,
			AVS_BURSTCOUNT_W          => 1,
			SUPPRESS_0_BYTEEN_CMD     => 1,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                        --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                 --       clk_reset.reset
			m0_address              => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_source0_ready,                                                                    --              cp.ready
			cp_valid                => burst_adapter_source0_valid,                                                                    --                .valid
			cp_data                 => burst_adapter_source0_data,                                                                     --                .data
			cp_startofpacket        => burst_adapter_source0_startofpacket,                                                            --                .startofpacket
			cp_endofpacket          => burst_adapter_source0_endofpacket,                                                              --                .endofpacket
			cp_channel              => burst_adapter_source0_channel,                                                                  --                .channel
			rf_sink_ready           => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                           --     (terminated)
			m0_writeresponserequest => open,                                                                                           --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                             --     (terminated)
		);

	lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 73,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                                        --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                 -- clk_reset.reset
			in_data           => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                           -- (terminated)
			csr_read          => '0',                                                                                            -- (terminated)
			csr_write         => '0',                                                                                            -- (terminated)
			csr_readdata      => open,                                                                                           -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                             -- (terminated)
			almost_full_data  => open,                                                                                           -- (terminated)
			almost_empty_data => open,                                                                                           -- (terminated)
			in_empty          => '0',                                                                                            -- (terminated)
			out_empty         => open,                                                                                           -- (terminated)
			in_error          => '0',                                                                                            -- (terminated)
			out_error         => open,                                                                                           -- (terminated)
			in_channel        => '0',                                                                                            -- (terminated)
			out_channel       => open                                                                                            -- (terminated)
		);

	addr_router : component lcd_addr_router
		port map (
			sink_ready         => master_0_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => master_0_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => master_0_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => master_0_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => master_0_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                     --       clk.clk
			reset              => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			src_ready          => addr_router_src_ready,                                                       --       src.ready
			src_valid          => addr_router_src_valid,                                                       --          .valid
			src_data           => addr_router_src_data,                                                        --          .data
			src_channel        => addr_router_src_channel,                                                     --          .channel
			src_startofpacket  => addr_router_src_startofpacket,                                               --          .startofpacket
			src_endofpacket    => addr_router_src_endofpacket                                                  --          .endofpacket
		);

	id_router : component lcd_id_router
		port map (
			sink_ready         => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => lcd_driver_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                              --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                       -- clk_reset.reset
			src_ready          => id_router_src_ready,                                                                  --       src.ready
			src_valid          => id_router_src_valid,                                                                  --          .valid
			src_data           => id_router_src_data,                                                                   --          .data
			src_channel        => id_router_src_channel,                                                                --          .channel
			src_startofpacket  => id_router_src_startofpacket,                                                          --          .startofpacket
			src_endofpacket    => id_router_src_endofpacket                                                             --          .endofpacket
		);

	burst_adapter : component altera_merlin_burst_adapter
		generic map (
			PKT_ADDR_H                => 40,
			PKT_ADDR_L                => 9,
			PKT_BEGIN_BURST           => 58,
			PKT_BYTE_CNT_H            => 49,
			PKT_BYTE_CNT_L            => 47,
			PKT_BYTEEN_H              => 8,
			PKT_BYTEEN_L              => 8,
			PKT_BURST_SIZE_H          => 53,
			PKT_BURST_SIZE_L          => 51,
			PKT_BURST_TYPE_H          => 55,
			PKT_BURST_TYPE_L          => 54,
			PKT_BURSTWRAP_H           => 50,
			PKT_BURSTWRAP_L           => 50,
			PKT_TRANS_COMPRESSED_READ => 41,
			PKT_TRANS_WRITE           => 43,
			PKT_TRANS_READ            => 44,
			OUT_NARROW_SIZE           => 0,
			IN_NARROW_SIZE            => 0,
			OUT_FIXED                 => 0,
			OUT_COMPLETE_WRAP         => 0,
			ST_DATA_W                 => 72,
			ST_CHANNEL_W              => 1,
			OUT_BYTE_CNT_H            => 47,
			OUT_BURSTWRAP_H           => 50,
			COMPRESSED_READ_SUPPORT   => 0,
			BYTEENABLE_SYNTHESIS      => 1,
			PIPE_INPUTS               => 0,
			NO_WRAP_SUPPORT           => 0,
			BURSTWRAP_CONST_MASK      => 1,
			BURSTWRAP_CONST_VALUE     => 1
		)
		port map (
			clk                   => clk_clk,                             --       cr0.clk
			reset                 => rst_controller_reset_out_reset,      -- cr0_reset.reset
			sink0_valid           => width_adapter_src_valid,             --     sink0.valid
			sink0_data            => width_adapter_src_data,              --          .data
			sink0_channel         => width_adapter_src_channel,           --          .channel
			sink0_startofpacket   => width_adapter_src_startofpacket,     --          .startofpacket
			sink0_endofpacket     => width_adapter_src_endofpacket,       --          .endofpacket
			sink0_ready           => width_adapter_src_ready,             --          .ready
			source0_valid         => burst_adapter_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_source0_data,          --          .data
			source0_channel       => burst_adapter_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_source0_ready          --          .ready
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS        => 1,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk        => clk_clk,                        --       clk.clk
			reset_out  => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req  => open,                           -- (terminated)
			reset_in1  => '0',                            -- (terminated)
			reset_in2  => '0',                            -- (terminated)
			reset_in3  => '0',                            -- (terminated)
			reset_in4  => '0',                            -- (terminated)
			reset_in5  => '0',                            -- (terminated)
			reset_in6  => '0',                            -- (terminated)
			reset_in7  => '0',                            -- (terminated)
			reset_in8  => '0',                            -- (terminated)
			reset_in9  => '0',                            -- (terminated)
			reset_in10 => '0',                            -- (terminated)
			reset_in11 => '0',                            -- (terminated)
			reset_in12 => '0',                            -- (terminated)
			reset_in13 => '0',                            -- (terminated)
			reset_in14 => '0',                            -- (terminated)
			reset_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS        => 1,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => lcd_clk_gen_0_reset_source_reset_ports_inv, -- reset_in0.reset
			clk        => clk_clk,                                    --       clk.clk
			reset_out  => rst_controller_001_reset_out_reset,         -- reset_out.reset
			reset_req  => open,                                       -- (terminated)
			reset_in1  => '0',                                        -- (terminated)
			reset_in2  => '0',                                        -- (terminated)
			reset_in3  => '0',                                        -- (terminated)
			reset_in4  => '0',                                        -- (terminated)
			reset_in5  => '0',                                        -- (terminated)
			reset_in6  => '0',                                        -- (terminated)
			reset_in7  => '0',                                        -- (terminated)
			reset_in8  => '0',                                        -- (terminated)
			reset_in9  => '0',                                        -- (terminated)
			reset_in10 => '0',                                        -- (terminated)
			reset_in11 => '0',                                        -- (terminated)
			reset_in12 => '0',                                        -- (terminated)
			reset_in13 => '0',                                        -- (terminated)
			reset_in14 => '0',                                        -- (terminated)
			reset_in15 => '0'                                         -- (terminated)
		);

	cmd_xbar_demux : component lcd_cmd_xbar_demux
		port map (
			clk                => clk_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,    -- clk_reset.reset
			sink_ready         => addr_router_src_ready,             --      sink.ready
			sink_channel       => addr_router_src_channel,           --          .channel
			sink_data          => addr_router_src_data,              --          .data
			sink_startofpacket => addr_router_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux : component lcd_cmd_xbar_demux
		port map (
			clk                => clk_clk,                             --       clk.clk
			reset              => rst_controller_reset_out_reset,      -- clk_reset.reset
			sink_ready         => width_adapter_001_src_ready,         --      sink.ready
			sink_channel       => width_adapter_001_src_channel,       --          .channel
			sink_data          => width_adapter_001_src_data,          --          .data
			sink_startofpacket => width_adapter_001_src_startofpacket, --          .startofpacket
			sink_endofpacket   => width_adapter_001_src_endofpacket,   --          .endofpacket
			sink_valid(0)      => width_adapter_001_src_valid,         --          .valid
			src0_ready         => rsp_xbar_demux_src0_ready,           --      src0.ready
			src0_valid         => rsp_xbar_demux_src0_valid,           --          .valid
			src0_data          => rsp_xbar_demux_src0_data,            --          .data
			src0_channel       => rsp_xbar_demux_src0_channel,         --          .channel
			src0_startofpacket => rsp_xbar_demux_src0_startofpacket,   --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_src0_endofpacket      --          .endofpacket
		);

	width_adapter : component lcd_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 67,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 76,
			IN_PKT_BYTE_CNT_L             => 74,
			IN_PKT_TRANS_COMPRESSED_READ  => 68,
			IN_PKT_BURSTWRAP_H            => 77,
			IN_PKT_BURSTWRAP_L            => 77,
			IN_PKT_BURST_SIZE_H           => 80,
			IN_PKT_BURST_SIZE_L           => 78,
			IN_PKT_RESPONSE_STATUS_H      => 98,
			IN_PKT_RESPONSE_STATUS_L      => 97,
			IN_PKT_TRANS_EXCLUSIVE        => 73,
			IN_PKT_BURST_TYPE_H           => 82,
			IN_PKT_BURST_TYPE_L           => 81,
			IN_ST_DATA_W                  => 99,
			OUT_PKT_ADDR_H                => 40,
			OUT_PKT_ADDR_L                => 9,
			OUT_PKT_DATA_H                => 7,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 8,
			OUT_PKT_BYTEEN_L              => 8,
			OUT_PKT_BYTE_CNT_H            => 49,
			OUT_PKT_BYTE_CNT_L            => 47,
			OUT_PKT_TRANS_COMPRESSED_READ => 41,
			OUT_PKT_BURST_SIZE_H          => 53,
			OUT_PKT_BURST_SIZE_L          => 51,
			OUT_PKT_RESPONSE_STATUS_H     => 71,
			OUT_PKT_RESPONSE_STATUS_L     => 70,
			OUT_PKT_TRANS_EXCLUSIVE       => 46,
			OUT_PKT_BURST_TYPE_H          => 55,
			OUT_PKT_BURST_TYPE_L          => 54,
			OUT_ST_DATA_W                 => 72,
			ST_CHANNEL_W                  => 1,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => clk_clk,                           --       clk.clk
			reset                => rst_controller_reset_out_reset,    -- clk_reset.reset
			in_valid             => cmd_xbar_demux_src0_valid,         --      sink.valid
			in_channel           => cmd_xbar_demux_src0_channel,       --          .channel
			in_startofpacket     => cmd_xbar_demux_src0_startofpacket, --          .startofpacket
			in_endofpacket       => cmd_xbar_demux_src0_endofpacket,   --          .endofpacket
			in_ready             => cmd_xbar_demux_src0_ready,         --          .ready
			in_data              => cmd_xbar_demux_src0_data,          --          .data
			out_endofpacket      => width_adapter_src_endofpacket,     --       src.endofpacket
			out_data             => width_adapter_src_data,            --          .data
			out_channel          => width_adapter_src_channel,         --          .channel
			out_valid            => width_adapter_src_valid,           --          .valid
			out_ready            => width_adapter_src_ready,           --          .ready
			out_startofpacket    => width_adapter_src_startofpacket,   --          .startofpacket
			in_command_size_data => "000"                              -- (terminated)
		);

	width_adapter_001 : component lcd_width_adapter_001
		generic map (
			IN_PKT_ADDR_H                 => 40,
			IN_PKT_ADDR_L                 => 9,
			IN_PKT_DATA_H                 => 7,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 8,
			IN_PKT_BYTEEN_L               => 8,
			IN_PKT_BYTE_CNT_H             => 49,
			IN_PKT_BYTE_CNT_L             => 47,
			IN_PKT_TRANS_COMPRESSED_READ  => 41,
			IN_PKT_BURSTWRAP_H            => 50,
			IN_PKT_BURSTWRAP_L            => 50,
			IN_PKT_BURST_SIZE_H           => 53,
			IN_PKT_BURST_SIZE_L           => 51,
			IN_PKT_RESPONSE_STATUS_H      => 71,
			IN_PKT_RESPONSE_STATUS_L      => 70,
			IN_PKT_TRANS_EXCLUSIVE        => 46,
			IN_PKT_BURST_TYPE_H           => 55,
			IN_PKT_BURST_TYPE_L           => 54,
			IN_ST_DATA_W                  => 72,
			OUT_PKT_ADDR_H                => 67,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 76,
			OUT_PKT_BYTE_CNT_L            => 74,
			OUT_PKT_TRANS_COMPRESSED_READ => 68,
			OUT_PKT_BURST_SIZE_H          => 80,
			OUT_PKT_BURST_SIZE_L          => 78,
			OUT_PKT_RESPONSE_STATUS_H     => 98,
			OUT_PKT_RESPONSE_STATUS_L     => 97,
			OUT_PKT_TRANS_EXCLUSIVE       => 73,
			OUT_PKT_BURST_TYPE_H          => 82,
			OUT_PKT_BURST_TYPE_L          => 81,
			OUT_ST_DATA_W                 => 99,
			ST_CHANNEL_W                  => 1,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => clk_clk,                             --       clk.clk
			reset                => rst_controller_reset_out_reset,      -- clk_reset.reset
			in_valid             => id_router_src_valid,                 --      sink.valid
			in_channel           => id_router_src_channel,               --          .channel
			in_startofpacket     => id_router_src_startofpacket,         --          .startofpacket
			in_endofpacket       => id_router_src_endofpacket,           --          .endofpacket
			in_ready             => id_router_src_ready,                 --          .ready
			in_data              => id_router_src_data,                  --          .data
			out_endofpacket      => width_adapter_001_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_001_src_data,          --          .data
			out_channel          => width_adapter_001_src_channel,       --          .channel
			out_valid            => width_adapter_001_src_valid,         --          .valid
			out_ready            => width_adapter_001_src_ready,         --          .ready
			out_startofpacket    => width_adapter_001_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	lcd_clk_gen_0_reset_source_reset_ports_inv <= not lcd_clk_gen_0_reset_source_reset;

end architecture rtl; -- of lcd
