library ieee;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity UART_LCD_Avalon_Master is
port (

);

end UART_LCD_Avalon_Master;

architecture struct of UART_LCD_Avalon_Master is

begin

end struct;